
module uart ( sys_clk, sys_rst_l, uart_XMIT_dataH, xmitH, xmit_dataH, 
        xmit_doneH, uart_REC_dataH, rec_dataH, rec_readyH, test_mode, test_se, 
        test_si, test_so );
  input [7:0] xmit_dataH;
  output [7:0] rec_dataH;
  input sys_clk, sys_rst_l, xmitH, uart_REC_dataH, test_mode, test_se, test_si;
  output uart_XMIT_dataH, xmit_doneH, rec_readyH, test_so;
  wire   iXMIT_xmit_doneInH, iXMIT_next_state_0_, iXMIT_next_state_1_,
         iXMIT_next_state_2_, iXMIT_state_0_, iXMIT_state_2_,
         iXMIT_bitCountH_0_, iXMIT_bitCountH_1_, iXMIT_bitCountH_2_,
         iXMIT_bitCountH_3_, iXMIT_N29, iXMIT_N28, iXMIT_N27, iXMIT_N26,
         iXMIT_bitCell_cntrH_0_, iXMIT_bitCell_cntrH_1_,
         iXMIT_bitCell_cntrH_2_, iXMIT_bitCell_cntrH_3_,
         iXMIT_xmit_ShiftRegH_1_, iXMIT_xmit_ShiftRegH_2_,
         iXMIT_xmit_ShiftRegH_3_, iXMIT_xmit_ShiftRegH_4_,
         iXMIT_xmit_ShiftRegH_5_, iXMIT_xmit_ShiftRegH_6_,
         iXMIT_xmit_ShiftRegH_7_, iRECEIVER_rec_readyInH,
         iRECEIVER_next_state_0_, iRECEIVER_next_state_1_,
         iRECEIVER_next_state_2_, iRECEIVER_state_0_, iRECEIVER_state_1_,
         iRECEIVER_state_2_, iRECEIVER_recd_bitCntrH_0_,
         iRECEIVER_recd_bitCntrH_1_, iRECEIVER_recd_bitCntrH_2_,
         iRECEIVER_recd_bitCntrH_3_, iRECEIVER_N23, iRECEIVER_N22,
         iRECEIVER_N21, iRECEIVER_N20, iRECEIVER_bitCell_cntrH_0_,
         iRECEIVER_bitCell_cntrH_1_, iRECEIVER_bitCell_cntrH_2_,
         iRECEIVER_bitCell_cntrH_3_, iRECEIVER_rec_datSyncH,
         iRECEIVER_rec_datH, n100, n103, n106, n109, n116, n123, n130, n137,
         n144, n151, n158, n165, n190, n193, n196, n199, n202, n205, n208,
         n211, n214, n217, n220, n223, n238, n239, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, \test_point/TM , n281,
         xmit_doneH_temp, rec_dataH_rec_0_temp, iXMIT_state_1_temp, n401, n94,
         n93, n92, n91, n9, n89, n88, n87, n86, n85, n84, n83, n82, n81, n80,
         n8, n79, n77, n75, n74, n73, n72, n71, n7, n69, n68, n67, n66, n65,
         n64, n63, n62, n61, n60, n58, n57, n56, n55, n54, n53, n52, n51, n50,
         n49, n48, n47, n46, n45, n44, n43, n42, n41, n39, n37, n35, n33, n31,
         n3, n29, n28, n275, n274, n273, n272, n271, n270, n27, n269, n268,
         n26, n25, n24, n23, n22, n21, n20, n2, n19, n18, n17, n15, n12, n11,
         n10, iXMIT_xmit_CTRL, iXMIT_state_1_, iXMIT_N_CTRL_2_,
         iXMIT_N_CTRL_1_, iXMIT_N46, iXMIT_N45, iXMIT_N44, iXMIT_N25,
         iXMIT_N24, iXMIT_N23, iXMIT_CRTL, iRECEIVER_state_CTRL,
         iRECEIVER_bitCell_CTRL, iRECEIVER_N_CTRL_2_, iRECEIVER_N_CTRL_1_,
         iRECEIVER_N28, iRECEIVER_N27, iRECEIVER_N26, iRECEIVER_N19,
         iRECEIVER_N18, iRECEIVER_N17, iRECEIVER_CTRL, iCTRL,
         \test_point/DOUT , n371, n370, n1, n6, n118, n119, n120, n121, n122,
         n124, n125, n126, n127, n128, n129, n131, n132, n133, n134, n135,
         n136, n138, n139, n140, n141, n142, n143, n145, n146, n147, n148,
         n149, n150, n152, n153, n154, n155, n156, n157, n159, n160, n161,
         n162, n163, n164, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182;
  wire   [7:0] rec_dataH_rec;
  wire   [7:0] rec_dataH_temp;
  assign \test_point/TM  = test_mode;
  assign test_so = rec_dataH_temp[7];

  AND2X4 U305 ( .IN1(iCTRL), .IN2(iXMIT_state_1_temp), .Q(iXMIT_state_1_) );
  AND2X4 U303 ( .IN1(iCTRL), .IN2(xmit_doneH_temp), .Q(xmit_doneH) );
  ISOLORX8 U302 ( .D(iXMIT_CRTL), .ISO(iRECEIVER_CTRL), .Q(iCTRL) );
  OR4X4 U301 ( .IN1(iRECEIVER_state_CTRL), .IN2(iRECEIVER_N_CTRL_1_), .IN3(
        iRECEIVER_N_CTRL_2_), .IN4(iRECEIVER_bitCell_CTRL), .Q(iRECEIVER_CTRL)
         );
  NAND4X1 U300 ( .IN1(iRECEIVER_N18), .IN2(iRECEIVER_N17), .IN3(
        iRECEIVER_bitCell_cntrH_0_), .IN4(iRECEIVER_bitCell_cntrH_1_), .QN(
        iRECEIVER_bitCell_CTRL) );
  NAND4X1 U299 ( .IN1(iRECEIVER_N22), .IN2(iRECEIVER_N21), .IN3(iRECEIVER_N20), 
        .IN4(iRECEIVER_N19), .QN(iRECEIVER_N_CTRL_2_) );
  NAND4X1 U298 ( .IN1(iRECEIVER_N28), .IN2(iRECEIVER_N27), .IN3(iRECEIVER_N26), 
        .IN4(iRECEIVER_N23), .QN(iRECEIVER_N_CTRL_1_) );
  NAND4X1 U297 ( .IN1(iRECEIVER_next_state_2_), .IN2(iRECEIVER_state_0_), 
        .IN3(iRECEIVER_state_1_), .IN4(iRECEIVER_state_2_), .QN(
        iRECEIVER_state_CTRL) );
  OR4X4 U296 ( .IN1(1'b0), .IN2(iXMIT_N_CTRL_1_), .IN3(iXMIT_N_CTRL_2_), .IN4(
        iXMIT_xmit_CTRL), .Q(iXMIT_CRTL) );
  NAND4X1 U295 ( .IN1(iXMIT_N24), .IN2(iXMIT_xmit_ShiftRegH_7_), .IN3(
        iXMIT_xmit_ShiftRegH_6_), .IN4(iXMIT_xmit_ShiftRegH_5_), .QN(
        iXMIT_xmit_CTRL) );
  NAND4X1 U294 ( .IN1(iXMIT_N28), .IN2(iXMIT_N27), .IN3(iXMIT_N26), .IN4(
        iXMIT_N25), .QN(iXMIT_N_CTRL_2_) );
  NAND4X1 U293 ( .IN1(n401), .IN2(n239), .IN3(n242), .IN4(n246), .QN(
        iXMIT_N_CTRL_1_) );
  XOR2X2 U230 ( .IN1(iRECEIVER_recd_bitCntrH_3_), .IN2(n275), .Q(iRECEIVER_N28) );
  NOR2X4 U229 ( .IN1(n274), .IN2(n250), .QN(n275) );
  XOR2X2 U228 ( .IN1(n250), .IN2(n274), .Q(iRECEIVER_N27) );
  XOR2X2 U227 ( .IN1(iRECEIVER_recd_bitCntrH_1_), .IN2(
        iRECEIVER_recd_bitCntrH_0_), .Q(iRECEIVER_N26) );
  XOR2X2 U226 ( .IN1(iRECEIVER_bitCell_cntrH_3_), .IN2(n273), .Q(iRECEIVER_N19) );
  NOR2X4 U225 ( .IN1(n272), .IN2(n249), .QN(n273) );
  XOR2X2 U224 ( .IN1(n249), .IN2(n272), .Q(iRECEIVER_N18) );
  XOR2X2 U223 ( .IN1(iRECEIVER_bitCell_cntrH_1_), .IN2(
        iRECEIVER_bitCell_cntrH_0_), .Q(iRECEIVER_N17) );
  XOR2X2 U222 ( .IN1(iXMIT_bitCountH_3_), .IN2(n271), .Q(iXMIT_N46) );
  NOR2X4 U221 ( .IN1(n270), .IN2(n247), .QN(n271) );
  XOR2X2 U220 ( .IN1(n247), .IN2(n270), .Q(iXMIT_N45) );
  XOR2X2 U219 ( .IN1(iXMIT_bitCountH_1_), .IN2(iXMIT_bitCountH_0_), .Q(
        iXMIT_N44) );
  XOR2X2 U218 ( .IN1(iXMIT_bitCell_cntrH_3_), .IN2(n269), .Q(iXMIT_N25) );
  NOR2X4 U217 ( .IN1(n268), .IN2(n251), .QN(n269) );
  XOR2X2 U216 ( .IN1(n251), .IN2(n268), .Q(iXMIT_N24) );
  XOR2X2 U215 ( .IN1(iXMIT_bitCell_cntrH_1_), .IN2(iXMIT_bitCell_cntrH_0_), 
        .Q(iXMIT_N23) );
  INVX32 U214 ( .INP(n64), .ZN(n28) );
  NAND2X4 U213 ( .IN1(n55), .IN2(n56), .QN(iXMIT_xmit_doneInH) );
  NAND2X4 U212 ( .IN1(iRECEIVER_bitCell_cntrH_1_), .IN2(
        iRECEIVER_bitCell_cntrH_0_), .QN(n272) );
  NAND2X4 U211 ( .IN1(iXMIT_bitCell_cntrH_1_), .IN2(iXMIT_bitCell_cntrH_0_), 
        .QN(n268) );
  NAND2X4 U210 ( .IN1(iRECEIVER_recd_bitCntrH_1_), .IN2(
        iRECEIVER_recd_bitCntrH_0_), .QN(n274) );
  NAND2X4 U209 ( .IN1(n61), .IN2(n69), .QN(n53) );
  NAND2X4 U208 ( .IN1(iXMIT_bitCountH_1_), .IN2(iXMIT_bitCountH_0_), .QN(n270)
         );
  NAND2X4 U207 ( .IN1(n63), .IN2(n44), .QN(iXMIT_next_state_1_) );
  NAND2X4 U206 ( .IN1(xmit_dataH[7]), .IN2(n26), .QN(n43) );
  NAND2X4 U205 ( .IN1(n42), .IN2(n43), .QN(n211) );
  NAND2X4 U204 ( .IN1(n67), .IN2(n68), .QN(iXMIT_next_state_0_) );
  INVX32 U202 ( .INP(n8), .ZN(n18) );
  NAND2X4 U201 ( .IN1(n80), .IN2(n91), .QN(n83) );
  NAND4X1 U138 ( .IN1(iRECEIVER_bitCell_cntrH_3_), .IN2(
        iRECEIVER_bitCell_cntrH_2_), .IN3(iRECEIVER_bitCell_cntrH_1_), .IN4(
        n255), .QN(n91) );
  INVX32 U137 ( .INP(n91), .ZN(n79) );
  AOI21X2 U135 ( .IN1(n79), .IN2(iRECEIVER_state_0_), .IN3(n241), .QN(n93) );
  NAND4X1 U132 ( .IN1(iRECEIVER_bitCell_cntrH_2_), .IN2(n255), .IN3(n244), 
        .IN4(n256), .QN(n85) );
  INVX32 U131 ( .INP(n85), .ZN(n88) );
  AOI21X2 U129 ( .IN1(n88), .IN2(n245), .IN3(iRECEIVER_state_2_), .QN(n94) );
  AND2X4 U128 ( .IN1(n93), .IN2(n94), .Q(n92) );
  AND2X4 U127 ( .IN1(n255), .IN2(n92), .Q(iRECEIVER_N20) );
  AND2X4 U126 ( .IN1(iRECEIVER_N17), .IN2(n92), .Q(iRECEIVER_N21) );
  AND2X4 U125 ( .IN1(iRECEIVER_N18), .IN2(n92), .Q(iRECEIVER_N22) );
  AND2X4 U124 ( .IN1(iRECEIVER_N19), .IN2(n92), .Q(iRECEIVER_N23) );
  NOR2X4 U123 ( .IN1(n241), .IN2(n245), .QN(n80) );
  NOR2X4 U120 ( .IN1(iRECEIVER_recd_bitCntrH_2_), .IN2(
        iRECEIVER_recd_bitCntrH_1_), .QN(n89) );
  NAND4X1 U118 ( .IN1(n80), .IN2(iRECEIVER_recd_bitCntrH_3_), .IN3(n89), .IN4(
        n243), .QN(n86) );
  AOI22X2 U117 ( .IN1(n88), .IN2(iRECEIVER_state_1_), .IN3(iRECEIVER_rec_datH), 
        .IN4(n241), .QN(n87) );
  NAND4X1 U116 ( .IN1(n83), .IN2(n238), .IN3(n86), .IN4(n87), .QN(
        iRECEIVER_next_state_0_) );
  AOI21X2 U114 ( .IN1(iRECEIVER_state_1_), .IN2(n85), .IN3(n248), .QN(n84) );
  ISOLORX8 U113 ( .D(iRECEIVER_state_0_), .ISO(n84), .Q(n81) );
  NAND3X4 U112 ( .IN1(n241), .IN2(n238), .IN3(n248), .QN(n82) );
  NOR2X4 U111 ( .IN1(n238), .IN2(iRECEIVER_state_0_), .QN(n8) );
  NAND4X1 U109 ( .IN1(n81), .IN2(n82), .IN3(n18), .IN4(n83), .QN(
        iRECEIVER_next_state_1_) );
  AND2X4 U108 ( .IN1(n79), .IN2(n80), .Q(iRECEIVER_next_state_2_) );
  NAND3X4 U107 ( .IN1(n241), .IN2(n238), .IN3(iRECEIVER_rec_datH), .QN(n77) );
  OAI21X2 U106 ( .IN1(n238), .IN2(n245), .IN3(n77), .QN(iRECEIVER_rec_readyInH) );
  NAND3X4 U102 ( .IN1(iXMIT_bitCell_cntrH_2_), .IN2(iXMIT_bitCell_cntrH_1_), 
        .IN3(iXMIT_bitCell_cntrH_3_), .QN(n75) );
  NOR2X4 U101 ( .IN1(n254), .IN2(n75), .QN(n57) );
  NOR2X4 U100 ( .IN1(n242), .IN2(n57), .QN(n62) );
  INVX32 U99 ( .INP(n62), .ZN(n72) );
  NOR2X4 U97 ( .IN1(n246), .IN2(iXMIT_state_0_), .QN(n66) );
  INVX32 U96 ( .INP(n57), .ZN(n74) );
  NOR2X4 U95 ( .IN1(n246), .IN2(n239), .QN(n54) );
  NOR2X4 U94 ( .IN1(n75), .IN2(iXMIT_bitCell_cntrH_0_), .QN(n61) );
  INVX32 U93 ( .INP(n61), .ZN(n65) );
  AOI22X2 U92 ( .IN1(n66), .IN2(n74), .IN3(n54), .IN4(n65), .QN(n73) );
  OAI21X2 U91 ( .IN1(n239), .IN2(n72), .IN3(n73), .QN(n71) );
  AND2X4 U90 ( .IN1(n254), .IN2(n71), .Q(iXMIT_N26) );
  AND2X4 U89 ( .IN1(iXMIT_N23), .IN2(n71), .Q(iXMIT_N27) );
  AND2X4 U88 ( .IN1(iXMIT_N24), .IN2(n71), .Q(iXMIT_N28) );
  AND2X4 U87 ( .IN1(iXMIT_N25), .IN2(n71), .Q(iXMIT_N29) );
  OR4X4 U85 ( .IN1(n253), .IN2(iXMIT_bitCountH_0_), .IN3(iXMIT_bitCountH_1_), 
        .IN4(iXMIT_bitCountH_2_), .Q(n69) );
  AOI22X2 U83 ( .IN1(n54), .IN2(n53), .IN3(iXMIT_state_2_), .IN4(n239), .QN(
        n67) );
  AOI21X2 U82 ( .IN1(n66), .IN2(n57), .IN3(n62), .QN(n68) );
  AOI21X2 U80 ( .IN1(iXMIT_state_1_temp), .IN2(n65), .IN3(n66), .QN(n63) );
  NAND3X4 U79 ( .IN1(n246), .IN2(n242), .IN3(xmitH), .QN(n64) );
  AOI21X2 U77 ( .IN1(n239), .IN2(iXMIT_state_2_), .IN3(n28), .QN(n44) );
  AOI22X2 U75 ( .IN1(n54), .IN2(n61), .IN3(n62), .IN4(iXMIT_state_0_), .QN(n60) );
  INVX32 U74 ( .INP(n60), .ZN(iXMIT_next_state_2_) );
  INVX32 U73 ( .INP(xmitH), .ZN(n58) );
  NAND3X4 U72 ( .IN1(n242), .IN2(n58), .IN3(n246), .QN(n55) );
  NAND3X4 U71 ( .IN1(iXMIT_state_2_), .IN2(iXMIT_state_0_), .IN3(n57), .QN(n56) );
  INVX32 U69 ( .INP(n55), .ZN(n51) );
  INVX32 U68 ( .INP(n54), .ZN(n52) );
  NOR2X4 U67 ( .IN1(n52), .IN2(n53), .QN(n47) );
  NOR2X4 U66 ( .IN1(n51), .IN2(n47), .QN(n46) );
  AOI22X2 U65 ( .IN1(iXMIT_bitCountH_0_), .IN2(n46), .IN3(n252), .IN4(n47), 
        .QN(n50) );
  INVX32 U64 ( .INP(n50), .ZN(n223) );
  AOI22X2 U63 ( .IN1(iXMIT_bitCountH_1_), .IN2(n46), .IN3(iXMIT_N44), .IN4(n47), .QN(n49) );
  INVX32 U62 ( .INP(n49), .ZN(n220) );
  AOI22X2 U61 ( .IN1(iXMIT_bitCountH_2_), .IN2(n46), .IN3(iXMIT_N45), .IN4(n47), .QN(n48) );
  INVX32 U60 ( .INP(n48), .ZN(n217) );
  AOI22X2 U59 ( .IN1(n46), .IN2(iXMIT_bitCountH_3_), .IN3(iXMIT_N46), .IN4(n47), .QN(n45) );
  INVX32 U58 ( .INP(n45), .ZN(n214) );
  NOR2X4 U57 ( .IN1(n44), .IN2(n28), .QN(n29) );
  AOI21X2 U56 ( .IN1(iXMIT_xmit_ShiftRegH_7_), .IN2(n44), .IN3(n29), .QN(n42)
         );
  INVX32 U55 ( .INP(n44), .ZN(n26) );
  AOI22X2 U51 ( .IN1(xmit_dataH[6]), .IN2(n28), .IN3(iXMIT_xmit_ShiftRegH_7_), 
        .IN4(n29), .QN(n41) );
  OAI21X2 U50 ( .IN1(n26), .IN2(n258), .IN3(n41), .QN(n208) );
  AOI22X2 U48 ( .IN1(xmit_dataH[5]), .IN2(n28), .IN3(iXMIT_xmit_ShiftRegH_6_), 
        .IN4(n29), .QN(n39) );
  OAI21X2 U47 ( .IN1(n26), .IN2(n259), .IN3(n39), .QN(n205) );
  AOI22X2 U45 ( .IN1(xmit_dataH[4]), .IN2(n28), .IN3(iXMIT_xmit_ShiftRegH_5_), 
        .IN4(n29), .QN(n37) );
  OAI21X2 U44 ( .IN1(n26), .IN2(n260), .IN3(n37), .QN(n202) );
  AOI22X2 U42 ( .IN1(xmit_dataH[3]), .IN2(n28), .IN3(iXMIT_xmit_ShiftRegH_4_), 
        .IN4(n29), .QN(n35) );
  OAI21X2 U41 ( .IN1(n26), .IN2(n261), .IN3(n35), .QN(n199) );
  AOI22X2 U39 ( .IN1(xmit_dataH[2]), .IN2(n28), .IN3(iXMIT_xmit_ShiftRegH_3_), 
        .IN4(n29), .QN(n33) );
  OAI21X2 U38 ( .IN1(n26), .IN2(n262), .IN3(n33), .QN(n196) );
  AOI22X2 U36 ( .IN1(xmit_dataH[1]), .IN2(n28), .IN3(iXMIT_xmit_ShiftRegH_2_), 
        .IN4(n29), .QN(n31) );
  OAI21X2 U35 ( .IN1(n263), .IN2(n26), .IN3(n31), .QN(n193) );
  AOI22X2 U33 ( .IN1(xmit_dataH[0]), .IN2(n28), .IN3(iXMIT_xmit_ShiftRegH_1_), 
        .IN4(n29), .QN(n27) );
  OAI21X2 U32 ( .IN1(n257), .IN2(n26), .IN3(n27), .QN(n190) );
  AOI22X2 U31 ( .IN1(iRECEIVER_rec_datH), .IN2(n8), .IN3(rec_dataH_rec[7]), 
        .IN4(n18), .QN(n25) );
  INVX32 U30 ( .INP(n25), .ZN(n165) );
  AOI22X2 U29 ( .IN1(rec_dataH_rec[7]), .IN2(n8), .IN3(rec_dataH_rec[6]), 
        .IN4(n18), .QN(n24) );
  INVX32 U28 ( .INP(n24), .ZN(n158) );
  AOI22X2 U27 ( .IN1(rec_dataH_rec[6]), .IN2(n8), .IN3(rec_dataH_rec[5]), 
        .IN4(n18), .QN(n23) );
  INVX32 U26 ( .INP(n23), .ZN(n151) );
  AOI22X2 U25 ( .IN1(rec_dataH_rec[5]), .IN2(n8), .IN3(rec_dataH_rec[4]), 
        .IN4(n18), .QN(n22) );
  INVX32 U24 ( .INP(n22), .ZN(n144) );
  AOI22X2 U23 ( .IN1(rec_dataH_rec[4]), .IN2(n8), .IN3(rec_dataH_rec[3]), 
        .IN4(n18), .QN(n21) );
  INVX32 U22 ( .INP(n21), .ZN(n137) );
  AOI22X2 U21 ( .IN1(rec_dataH_rec[3]), .IN2(n8), .IN3(rec_dataH_rec[2]), 
        .IN4(n18), .QN(n20) );
  INVX32 U20 ( .INP(n20), .ZN(n130) );
  AOI22X2 U19 ( .IN1(rec_dataH_rec[2]), .IN2(n8), .IN3(rec_dataH_rec[1]), 
        .IN4(n18), .QN(n19) );
  INVX32 U18 ( .INP(n19), .ZN(n123) );
  AOI22X2 U17 ( .IN1(rec_dataH_rec[1]), .IN2(n8), .IN3(rec_dataH_rec_0_temp), 
        .IN4(n18), .QN(n17) );
  INVX32 U16 ( .INP(n17), .ZN(n116) );
  OAI21X2 U15 ( .IN1(iRECEIVER_state_1_), .IN2(n248), .IN3(n238), .QN(n15) );
  OAI21X2 U14 ( .IN1(n238), .IN2(n245), .IN3(n15), .QN(n9) );
  AOI22X2 U13 ( .IN1(iRECEIVER_N28), .IN2(n8), .IN3(iRECEIVER_recd_bitCntrH_3_), .IN4(n9), .QN(n12) );
  INVX32 U12 ( .INP(n12), .ZN(n109) );
  AOI22X2 U11 ( .IN1(n243), .IN2(n8), .IN3(iRECEIVER_recd_bitCntrH_0_), .IN4(
        n9), .QN(n11) );
  INVX32 U10 ( .INP(n11), .ZN(n106) );
  AOI22X2 U9 ( .IN1(iRECEIVER_N26), .IN2(n8), .IN3(iRECEIVER_recd_bitCntrH_1_), 
        .IN4(n9), .QN(n10) );
  INVX32 U8 ( .INP(n10), .ZN(n103) );
  AOI22X2 U7 ( .IN1(iRECEIVER_N27), .IN2(n8), .IN3(iRECEIVER_recd_bitCntrH_2_), 
        .IN4(n9), .QN(n7) );
  INVX32 U6 ( .INP(n7), .ZN(n100) );
  AOI21X2 U5 ( .IN1(n242), .IN2(n239), .IN3(n257), .QN(n3) );
  AOI21X2 U4 ( .IN1(iXMIT_state_2_), .IN2(iXMIT_state_0_), .IN3(n3), .QN(n2)
         );
  OAI21X2 U3 ( .IN1(iXMIT_state_2_), .IN2(iXMIT_state_1_), .IN3(n2), .QN(
        uart_XMIT_dataH) );
  INVX32 U290 ( .INP(n370), .ZN(n371) );
  NAND2X4 U289 ( .IN1(1'b1), .IN2(\test_point/TM ), .QN(n370) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_2_ ( .D(n182), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_bitCell_cntrH_2_), .QN(n251) );
  DFFARX1 iXMIT_state_reg_0_ ( .D(n181), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_0_), .QN(n239) );
  DFFARX1 iXMIT_state_reg_2_ ( .D(n180), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_2_), .QN(n242) );
  DFFARX1 iXMIT_state_reg_1_ ( .D(n179), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        iXMIT_state_1_temp), .QN(n246) );
  DFFARX1 iXMIT_bitCountH_reg_0_ ( .D(n178), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iXMIT_bitCountH_0_), .QN(n252) );
  DFFARX1 iXMIT_bitCountH_reg_1_ ( .D(n177), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iXMIT_bitCountH_1_) );
  DFFARX1 iXMIT_bitCountH_reg_2_ ( .D(n176), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iXMIT_bitCountH_2_), .QN(n247) );
  DFFARX1 iXMIT_bitCountH_reg_3_ ( .D(n175), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iXMIT_bitCountH_3_), .QN(n253) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_7_ ( .D(n174), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_7_) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_6_ ( .D(n173), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_6_), .QN(n258) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_5_ ( .D(n172), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_5_), .QN(n259) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_4_ ( .D(n171), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_4_), .QN(n260) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_3_ ( .D(n170), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_3_), .QN(n261) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_2_ ( .D(n169), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_2_), .QN(n262) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_1_ ( .D(n168), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_xmit_ShiftRegH_1_), .QN(n263) );
  DFFARX1 iXMIT_xmit_doneH_reg ( .D(n167), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(xmit_doneH_temp) );
  DFFARX1 iRECEIVER_state_reg_1_ ( .D(n166), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_1_), .QN(n241) );
  DFFASX1 iRECEIVER_state_reg_0_ ( .D(n164), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_state_0_), .QN(n245) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_0_ ( .D(n163), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_0_), .QN(n255) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_1_ ( .D(n162), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_1_), .QN(n244) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_2_ ( .D(n161), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_2_), .QN(n249) );
  DFFARX1 iRECEIVER_bitCell_cntrH_reg_3_ ( .D(n160), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_bitCell_cntrH_3_), .QN(n256) );
  DFFARX1 iRECEIVER_state_reg_2_ ( .D(n159), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(iRECEIVER_state_2_), .QN(n238) );
  DFFARX1 iRECEIVER_rec_readyH_reg ( .D(n157), .CLK(sys_clk), .RSTB(sys_rst_l), 
        .Q(rec_readyH) );
  DFFARX1 iRECEIVER_par_dataH_reg_7_ ( .D(n156), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec[7]) );
  DFFARX1 rec_dataH_temp_reg_7_ ( .D(n155), .CLK(\test_point/DOUT ), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp[7]) );
  DFFARX1 rec_dataH_reg_7_ ( .D(n154), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH[7]) );
  DFFARX1 iRECEIVER_par_dataH_reg_6_ ( .D(n153), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec[6]) );
  DFFARX1 rec_dataH_temp_reg_6_ ( .D(n152), .CLK(\test_point/DOUT ), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp[6]) );
  DFFARX1 rec_dataH_reg_6_ ( .D(n150), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH[6]) );
  DFFARX1 iRECEIVER_par_dataH_reg_5_ ( .D(n149), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec[5]) );
  DFFARX1 rec_dataH_temp_reg_5_ ( .D(n148), .CLK(\test_point/DOUT ), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp[5]) );
  DFFARX1 rec_dataH_reg_5_ ( .D(n147), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH[5]) );
  DFFARX1 iRECEIVER_par_dataH_reg_4_ ( .D(n146), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec[4]) );
  DFFARX1 rec_dataH_temp_reg_4_ ( .D(n145), .CLK(\test_point/DOUT ), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp[4]) );
  DFFARX1 rec_dataH_reg_4_ ( .D(n143), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH[4]) );
  DFFARX1 iRECEIVER_par_dataH_reg_3_ ( .D(n142), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec[3]) );
  DFFARX1 rec_dataH_temp_reg_3_ ( .D(n141), .CLK(\test_point/DOUT ), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp[3]) );
  DFFARX1 rec_dataH_reg_3_ ( .D(n140), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH[3]) );
  DFFARX1 iRECEIVER_par_dataH_reg_2_ ( .D(n139), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec[2]) );
  DFFARX1 rec_dataH_temp_reg_2_ ( .D(n138), .CLK(\test_point/DOUT ), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp[2]) );
  DFFARX1 rec_dataH_reg_2_ ( .D(n136), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH[2]) );
  DFFARX1 iRECEIVER_par_dataH_reg_1_ ( .D(n135), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec[1]) );
  DFFARX1 rec_dataH_temp_reg_1_ ( .D(n134), .CLK(\test_point/DOUT ), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp[1]) );
  DFFARX1 rec_dataH_reg_1_ ( .D(n133), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH[1]) );
  DFFARX1 iRECEIVER_par_dataH_reg_0_ ( .D(n132), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(rec_dataH_rec_0_temp) );
  DFFARX1 rec_dataH_temp_reg_0_ ( .D(n131), .CLK(\test_point/DOUT ), .RSTB(
        sys_rst_l), .Q(rec_dataH_temp[0]) );
  DFFARX1 rec_dataH_reg_0_ ( .D(n129), .CLK(sys_clk), .RSTB(sys_rst_l), .Q(
        rec_dataH[0]) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_3_ ( .D(n128), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_recd_bitCntrH_3_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_0_ ( .D(n127), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_recd_bitCntrH_0_), .QN(n243) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_1_ ( .D(n126), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_recd_bitCntrH_1_) );
  DFFARX1 iRECEIVER_recd_bitCntrH_reg_2_ ( .D(n125), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iRECEIVER_recd_bitCntrH_2_), .QN(n250) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_3_ ( .D(n124), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_bitCell_cntrH_3_) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_0_ ( .D(n122), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_bitCell_cntrH_0_), .QN(n254) );
  DFFARX1 iXMIT_bitCell_cntrH_reg_1_ ( .D(n121), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(iXMIT_bitCell_cntrH_1_), .QN(n6) );
  DFFARX1 iXMIT_xmit_ShiftRegH_reg_0_ ( .D(n120), .CLK(sys_clk), .RSTB(
        sys_rst_l), .Q(n281), .QN(n257) );
  DFFASX1 iRECEIVER_rec_datSyncH_reg ( .D(n119), .CLK(sys_clk), .SETB(
        sys_rst_l), .Q(iRECEIVER_rec_datSyncH) );
  DFFASX1 iRECEIVER_rec_datH_reg ( .D(n118), .CLK(sys_clk), .SETB(sys_rst_l), 
        .Q(iRECEIVER_rec_datH), .QN(n248) );
  DFFARX1 iDatasend_reg_2_ ( .D(n182), .CLK(sys_clk), .RSTB(sys_rst_l), .QN(
        n401) );
  MUX21X2 U291 ( .IN1(rec_readyH), .IN2(sys_clk), .S(n371), .Q(
        \test_point/DOUT ) );
  MUX21X1 U1 ( .IN1(iRECEIVER_N22), .IN2(iRECEIVER_bitCell_cntrH_1_), .S(
        test_se), .Q(n161) );
  MUX21X1 U2 ( .IN1(iRECEIVER_N21), .IN2(iRECEIVER_bitCell_cntrH_0_), .S(
        test_se), .Q(n162) );
  MUX21X1 U34 ( .IN1(iRECEIVER_N20), .IN2(test_si), .S(test_se), .Q(n163) );
  MUX21X1 U37 ( .IN1(iRECEIVER_next_state_0_), .IN2(iRECEIVER_recd_bitCntrH_3_), .S(test_se), .Q(n164) );
  MUX21X1 U40 ( .IN1(iRECEIVER_next_state_1_), .IN2(iRECEIVER_state_0_), .S(
        test_se), .Q(n166) );
  MUX21X1 U43 ( .IN1(iXMIT_xmit_doneInH), .IN2(iXMIT_xmit_ShiftRegH_7_), .S(
        test_se), .Q(n167) );
  MUX21X1 U46 ( .IN1(n193), .IN2(n281), .S(test_se), .Q(n168) );
  MUX21X1 U49 ( .IN1(n196), .IN2(iXMIT_xmit_ShiftRegH_1_), .S(test_se), .Q(
        n169) );
  MUX21X1 U52 ( .IN1(n199), .IN2(iXMIT_xmit_ShiftRegH_2_), .S(test_se), .Q(
        n170) );
  MUX21X1 U53 ( .IN1(n202), .IN2(iXMIT_xmit_ShiftRegH_3_), .S(test_se), .Q(
        n171) );
  MUX21X1 U54 ( .IN1(n205), .IN2(iXMIT_xmit_ShiftRegH_4_), .S(test_se), .Q(
        n172) );
  MUX21X1 U70 ( .IN1(n208), .IN2(iXMIT_xmit_ShiftRegH_5_), .S(test_se), .Q(
        n173) );
  MUX21X1 U76 ( .IN1(n211), .IN2(iXMIT_xmit_ShiftRegH_6_), .S(test_se), .Q(
        n174) );
  MUX21X1 U78 ( .IN1(n214), .IN2(iXMIT_bitCountH_2_), .S(test_se), .Q(n175) );
  MUX21X1 U81 ( .IN1(n217), .IN2(iXMIT_bitCountH_1_), .S(test_se), .Q(n176) );
  MUX21X1 U84 ( .IN1(n220), .IN2(iXMIT_bitCountH_0_), .S(test_se), .Q(n177) );
  MUX21X1 U86 ( .IN1(n223), .IN2(iXMIT_bitCell_cntrH_3_), .S(test_se), .Q(n178) );
  MUX21X1 U98 ( .IN1(iXMIT_next_state_1_), .IN2(iXMIT_state_0_), .S(test_se), 
        .Q(n179) );
  MUX21X1 U103 ( .IN1(iXMIT_next_state_2_), .IN2(iXMIT_state_1_temp), .S(
        test_se), .Q(n180) );
  MUX21X1 U104 ( .IN1(iXMIT_next_state_0_), .IN2(iXMIT_bitCountH_3_), .S(
        test_se), .Q(n181) );
  MUX21X1 U105 ( .IN1(iRECEIVER_rec_datSyncH), .IN2(rec_dataH_rec[7]), .S(
        test_se), .Q(n118) );
  MUX21X1 U110 ( .IN1(uart_REC_dataH), .IN2(iRECEIVER_rec_datH), .S(test_se), 
        .Q(n119) );
  MUX21X1 U115 ( .IN1(n190), .IN2(iXMIT_state_2_), .S(test_se), .Q(n120) );
  MUX21X1 U119 ( .IN1(iXMIT_N27), .IN2(iXMIT_bitCell_cntrH_0_), .S(test_se), 
        .Q(n121) );
  MUX21X1 U121 ( .IN1(iXMIT_N26), .IN2(iRECEIVER_state_2_), .S(test_se), .Q(
        n122) );
  MUX21X1 U122 ( .IN1(iXMIT_N29), .IN2(iXMIT_bitCell_cntrH_2_), .S(test_se), 
        .Q(n124) );
  MUX21X1 U130 ( .IN1(n100), .IN2(iRECEIVER_recd_bitCntrH_1_), .S(test_se), 
        .Q(n125) );
  MUX21X1 U133 ( .IN1(n103), .IN2(iRECEIVER_recd_bitCntrH_0_), .S(test_se), 
        .Q(n126) );
  MUX21X1 U134 ( .IN1(n106), .IN2(rec_readyH), .S(test_se), .Q(n127) );
  MUX21X1 U136 ( .IN1(n109), .IN2(iRECEIVER_recd_bitCntrH_2_), .S(test_se), 
        .Q(n128) );
  MUX21X1 U139 ( .IN1(rec_dataH_temp[0]), .IN2(xmit_doneH_temp), .S(test_se), 
        .Q(n129) );
  MUX21X1 U140 ( .IN1(rec_dataH_rec_0_temp), .IN2(rec_dataH[7]), .S(test_se), 
        .Q(n131) );
  MUX21X1 U141 ( .IN1(n116), .IN2(iRECEIVER_bitCell_cntrH_3_), .S(test_se), 
        .Q(n132) );
  MUX21X1 U142 ( .IN1(rec_dataH_temp[1]), .IN2(rec_dataH[0]), .S(test_se), .Q(
        n133) );
  MUX21X1 U143 ( .IN1(rec_dataH_rec[1]), .IN2(rec_dataH_temp[0]), .S(test_se), 
        .Q(n134) );
  MUX21X1 U144 ( .IN1(n123), .IN2(rec_dataH_rec_0_temp), .S(test_se), .Q(n135)
         );
  MUX21X1 U145 ( .IN1(rec_dataH_temp[2]), .IN2(rec_dataH[1]), .S(test_se), .Q(
        n136) );
  MUX21X1 U146 ( .IN1(rec_dataH_rec[2]), .IN2(rec_dataH_temp[1]), .S(test_se), 
        .Q(n138) );
  MUX21X1 U147 ( .IN1(n130), .IN2(rec_dataH_rec[1]), .S(test_se), .Q(n139) );
  MUX21X1 U148 ( .IN1(rec_dataH_temp[3]), .IN2(rec_dataH[2]), .S(test_se), .Q(
        n140) );
  MUX21X1 U149 ( .IN1(rec_dataH_rec[3]), .IN2(rec_dataH_temp[2]), .S(test_se), 
        .Q(n141) );
  MUX21X1 U150 ( .IN1(n137), .IN2(rec_dataH_rec[2]), .S(test_se), .Q(n142) );
  MUX21X1 U151 ( .IN1(rec_dataH_temp[4]), .IN2(rec_dataH[3]), .S(test_se), .Q(
        n143) );
  MUX21X1 U152 ( .IN1(rec_dataH_rec[4]), .IN2(rec_dataH_temp[3]), .S(test_se), 
        .Q(n145) );
  MUX21X1 U153 ( .IN1(n144), .IN2(rec_dataH_rec[3]), .S(test_se), .Q(n146) );
  MUX21X1 U154 ( .IN1(rec_dataH_temp[5]), .IN2(rec_dataH[4]), .S(test_se), .Q(
        n147) );
  MUX21X1 U155 ( .IN1(rec_dataH_rec[5]), .IN2(rec_dataH_temp[4]), .S(test_se), 
        .Q(n148) );
  MUX21X1 U156 ( .IN1(n151), .IN2(rec_dataH_rec[4]), .S(test_se), .Q(n149) );
  MUX21X1 U157 ( .IN1(rec_dataH_temp[6]), .IN2(rec_dataH[5]), .S(test_se), .Q(
        n150) );
  MUX21X1 U158 ( .IN1(rec_dataH_rec[6]), .IN2(rec_dataH_temp[5]), .S(test_se), 
        .Q(n152) );
  MUX21X1 U159 ( .IN1(n158), .IN2(rec_dataH_rec[5]), .S(test_se), .Q(n153) );
  MUX21X1 U160 ( .IN1(rec_dataH_temp[7]), .IN2(rec_dataH[6]), .S(test_se), .Q(
        n154) );
  MUX21X1 U161 ( .IN1(rec_dataH_rec[7]), .IN2(rec_dataH_temp[6]), .S(test_se), 
        .Q(n155) );
  MUX21X1 U162 ( .IN1(n165), .IN2(rec_dataH_rec[6]), .S(test_se), .Q(n156) );
  MUX21X1 U163 ( .IN1(iRECEIVER_rec_readyInH), .IN2(iRECEIVER_rec_datSyncH), 
        .S(test_se), .Q(n157) );
  MUX21X1 U164 ( .IN1(iRECEIVER_next_state_2_), .IN2(iRECEIVER_state_1_), .S(
        test_se), .Q(n159) );
  MUX21X1 U165 ( .IN1(iRECEIVER_N23), .IN2(iRECEIVER_bitCell_cntrH_2_), .S(
        test_se), .Q(n160) );
  MUX21X1 U166 ( .IN1(iXMIT_N28), .IN2(n1), .S(test_se), .Q(n182) );
  INVX0 U167 ( .INP(n6), .ZN(n1) );
endmodule

